class fifo_driver extends uvm_driver #(fifo_sequence_items);
  
