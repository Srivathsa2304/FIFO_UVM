class fifo_sequencer extends uvm_sequencer#(fifo_sequence_items);
