class fifo_sequence extends uvm_sequence #();
